module mod_c();
endmodule
