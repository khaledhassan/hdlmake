module level0;
  //level1 g();
endmodule
