`include "notfount.vh"

module gate;
  wire w3;
endmodule
