import pkg::*;

module gate;
  wire w3;
endmodule
