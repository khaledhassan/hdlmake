package test_pkg is
  constant C_TEST_INT : integer := 5;
end package;

