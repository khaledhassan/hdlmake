module level2;
  level1 g();
endmodule
