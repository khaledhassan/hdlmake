`include "macros.v"

module gate;
  initial
   $display("hello");
endmodule
