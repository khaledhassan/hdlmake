package pkg;
  const int v = 5;
endpackage;
