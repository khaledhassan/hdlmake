module gate2(input i, output o);
  assign o = ~i;
endmodule
