module mod2;
  logic v;
endmodule;
