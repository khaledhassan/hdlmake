`define one 1
`define include(x) x^1

module gate;
  wire w3;
endmodule
