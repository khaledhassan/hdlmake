context testlib_context is
  library testlib;
  use testlib.test_pkg.all;
end context;
