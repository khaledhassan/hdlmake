module mod_b();
endmodule
