module gate;
  level2 g();
  level1 h();
endmodule
