

module gate3(input a);
endmodule
