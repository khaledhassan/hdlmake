module gate;
  wire `name(w3);
endmodule
