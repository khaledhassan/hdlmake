module level1;
  level0 g();
endmodule
