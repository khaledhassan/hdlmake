use work.all;

entity gate is
end;

architecture arch of gate is
begin
   assert false report msg;
end arch;
