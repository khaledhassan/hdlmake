package pkg is
  constant msg : string := "hello";
end;

