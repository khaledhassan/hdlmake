module unused;
endmodule
