`define nest(x) `nest(x)

module gate;
  wire `nest(w3);
endmodule
