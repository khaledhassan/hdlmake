module mod_a();
endmodule
